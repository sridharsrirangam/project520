module changeInYMat();
